`include "test_base.vh"
`include "test_ldi.vh"
`include "test_lds.vh"
`include "test_sts.vh"
`include "test_ldy.vh"
`include "test_mov.vh"
`include "test_add.vh"
`include "test_sub.vh"
`include "test_pop.vh"
`include "test_push.vh"
`include "test_brbs.vh"
`include "test_brcs.vh"
`include "test_rjmp.vh"
`include "test_rcall.vh"
`include "test_ret.vh"